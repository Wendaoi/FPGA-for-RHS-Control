// =============================================================================
// 模块名称: data_input_module
// 描述:    数据输入模块，负责从RHS芯片捕获原始数据并进行预处理
//          根据电极分组配置决定是否捕获特定电极的数据
// =============================================================================

`timescale 1ns/1ps

module data_input_module #(
    parameter DATA_WIDTH = 16,          // 数据宽度 (默认16位)
    parameter CHANNELS = 8,             // 通道数量 (默认8通道)
    parameter GROUPS = 10,              // 电极分组数量 (默认10组)
    parameter ELECTRODES_PER_GROUP = 8  // 每组电极数量 (默认每组8个电极)
) (
    // -------------------------------------------------------------------------
    // 系统时钟和复位信号
    // -------------------------------------------------------------------------
    input wire clk,                     // 系统时钟
    input wire reset,                   // 系统复位信号 (高电平有效)
    
    // -------------------------------------------------------------------------
    // RHS芯片数据输入接口
    // 从RHS2000系列芯片接收原始生物电信号数据
    // -------------------------------------------------------------------------
    input wire [DATA_WIDTH-1:0] rhs_data_in [0:CHANNELS-1],  // RHS芯片数据输入 (每个通道DATA_WIDTH位)
    input wire rhs_data_valid,                               // RHS数据有效信号
    
    // -------------------------------------------------------------------------
    // 电极分组控制接口
    // 用于配置电极分组和功能，决定哪些电极需要捕获数据
    // -------------------------------------------------------------------------
    // 电极分组映射表
    // group_map[组号][电极号] = 实际电极编号
    input wire [7:0] group_map [0:GROUPS-1][0:ELECTRODES_PER_GROUP-1],
    
    // 电极功能配置数组
    // 每组电极的功能配置：
    // 00: 收集电位信号
    // 01: 发送刺激
    // 10: 高阻态
    // 11: 保留
    input wire [1:0] electrode_function [0:GROUPS-1],
    
    // 当前操作的组号 (0-9)
    input wire [3:0] current_group,
    
    // -------------------------------------------------------------------------
    // 数据输出接口
    // 向下游模块输出经过预处理的数据
    // -------------------------------------------------------------------------
    output reg [DATA_WIDTH-1:0] processed_data [0:CHANNELS-1],  // 经过预处理的数据
    output reg data_out_valid,                                   // 数据输出有效信号
    
    // -------------------------------------------------------------------------
    // 控制接口
    // 控制数据捕获的启动和完成状态反馈
    // -------------------------------------------------------------------------
    input wire data_capture_en,         // 数据捕获使能信号
    output reg data_capture_done         // 数据捕获完成信号
);

// -------------------------------------------------------------------------
// 内部信号定义
// -------------------------------------------------------------------------

// 状态机状态寄存器
reg [2:0] state;                                    // 当前状态 (3位状态机)

// 数据缓冲区
reg [DATA_WIDTH-1:0] data_buffer [0:CHANNELS-1];    // 数据缓冲区，存储从RHS芯片捕获的原始数据
reg data_buffer_valid;                              // 数据缓冲区有效标志

// -------------------------------------------------------------------------
// 状态机定义 - 控制数据捕获和处理的时序
// -------------------------------------------------------------------------

localparam IDLE = 3'd0;        // 空闲状态：等待数据捕获使能
localparam CAPTURE = 3'd1;     // 捕获状态：从RHS芯片捕获数据
localparam PROCESS = 3'd2;     // 处理状态：对捕获的数据进行预处理
localparam OUTPUT = 3'd3;      // 输出状态：向下游模块输出处理后的数据

// -------------------------------------------------------------------------
// 主要状态机逻辑 - 控制数据捕获、处理和输出的完整流程
// -------------------------------------------------------------------------

always @(posedge clk or posedge reset) begin
    if (reset) begin
        // ---------------------------------------------------------------------
        // 复位状态下初始化所有信号和状态
        // ---------------------------------------------------------------------
        state <= IDLE;                          // 状态机复位到空闲状态
        data_buffer_valid <= 1'b0;              // 数据缓冲区有效标志清零
        data_out_valid <= 1'b0;                 // 数据输出有效标志清零
        data_capture_done <= 1'b0;              // 数据捕获完成标志清零
        
        // ---------------------------------------------------------------------
        // 初始化数据缓冲区和输出数组
        // ---------------------------------------------------------------------
        integer i;
        for (i = 0; i < CHANNELS; i = i + 1) begin
            data_buffer[i] <= {DATA_WIDTH{1'b0}};      // 数据缓冲区清零
            processed_data[i] <= {DATA_WIDTH{1'b0}};    // 处理后数据清零
        end
    end else begin
        case (state)
            // ---------------------------------------------------------------------
            // IDLE状态 - 空闲状态
            // 等待数据捕获使能信号和有效的RHS数据
            // ---------------------------------------------------------------------
            IDLE: begin
                data_buffer_valid <= 1'b0;              // 清除数据缓冲区有效标志
                data_out_valid <= 1'b0;                 // 清除数据输出有效标志
                data_capture_done <= 1'b0;              // 清除数据捕获完成标志
                
                // 检查是否满足数据捕获条件
                if (data_capture_en && rhs_data_valid) begin
                    state <= CAPTURE;                   // 满足条件时转到捕获状态
                end
                // 否则继续保持空闲状态
            end
            
            // ---------------------------------------------------------------------
            // CAPTURE状态 - 数据捕获状态
            // 从RHS芯片捕获原始数据，根据电极分组配置决定是否捕获特定电极数据
            // ---------------------------------------------------------------------
            CAPTURE: begin
                // 捕获RHS芯片数据
                integer i;
                for (i = 0; i < CHANNELS; i = i + 1) begin
                    // -----------------------------------------------------------------
                    // 检查当前通道是否属于当前操作的组
                    // 如果属于当前组且功能为发送刺激，则不捕获数据
                    // -----------------------------------------------------------------
                    reg is_current_group_electrode;
                    integer g, e;
                    is_current_group_electrode = 1'b0;
                    
                    // 检查当前电极是否属于当前组
                    for (g = 0; g < GROUPS; g = g + 1) begin
                        for (e = 0; e < ELECTRODES_PER_GROUP; e = e + 1) begin
                            // 如果当前电极编号等于通道i，且组号等于当前操作组，且功能为发送刺激
                            if (group_map[g][e] == i && g == current_group && electrode_function[g] == 2'b01) begin
                                is_current_group_electrode = 1'b1;  // 标记为当前组的刺激电极
                            end
                        end
                    end
                    
                    // -----------------------------------------------------------------
                    // 根据电极功能决定是否捕获数据
                    // -----------------------------------------------------------------
                    // 如果不是当前组的刺激电极，则捕获数据
                    if (!is_current_group_electrode) begin
                        data_buffer[i] <= rhs_data_in[i];          // 捕获RHS芯片数据
                    end else begin
                        // 对于当前组的刺激电极，设置为默认值（不捕获数据）
                        data_buffer[i] <= {DATA_WIDTH{1'b0}};      // 设置为零值
                    end
                end
                data_buffer_valid <= 1'b1;                         // 设置数据缓冲区有效标志
                state <= PROCESS;                                   // 转到处理状态
            end
            
            // ---------------------------------------------------------------------
            // PROCESS状态 - 数据处理状态
            // 对捕获的数据进行预处理（当前版本为直通处理）
            // ---------------------------------------------------------------------
            PROCESS: begin
                // 数据预处理（这里可以添加更多处理逻辑）
                integer i;
                for (i = 0; i < CHANNELS; i = i + 1) begin
                    processed_data[i] <= data_buffer[i];            // 直接复制缓冲区数据到输出
                end
                data_out_valid <= 1'b1;                             // 设置数据输出有效标志
                data_capture_done <= 1'b1;                          // 设置数据捕获完成标志
                state <= OUTPUT;                                    // 转到输出状态
            end
            
            // ---------------------------------------------------------------------
            // OUTPUT状态 - 数据输出状态
            // 保持输出状态直到上游模块消费数据
            // ---------------------------------------------------------------------
            OUTPUT: begin
                // 保持输出状态直到数据被消费
                if (!data_capture_en) begin
                    data_out_valid <= 1'b0;                         // 清除数据输出有效标志
                    data_capture_done <= 1'b0;                      // 清除数据捕获完成标志
                    state <= IDLE;                                  // 返回空闲状态
                end
                // 否则继续保持输出状态
            end
        endcase
    end
end

endmodule